module control (
	input [5:0] op,

	output reg memread, memwrite, alusrca, memtoreg, iord, regwrite, regdest,
	output pcen,
	output reg [1:0] pcsource, alusrcb, aluop,
	output reg [3:0] iwrite
);

	

endmodule;