module control (
	input [5:0] op,

	output out
);

endmodule;