module register_file (
	input [1:0] 	read_adr_a,
	input [1:0] 	read_adr_b,
	input [1:0] 	write_adr,
	input [47:0]	write_data,
	input 			write_en,

	output [47:0] 	reg_a,
	output [47:0] 	reg_b
);



endmodule